module craft_encrypt (
    input wire clk,
    input wire rst,
    input wire [63:0] plaintext,
    input wire [63:0] tweak,
    input wire [127:0] key,
    output wire done,
    output wire [63:0] ciphertext
);



endmodule  //craft_encrypt
