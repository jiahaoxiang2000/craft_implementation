module craft_state_register (
    input clk,
    input en
);

endmodule
